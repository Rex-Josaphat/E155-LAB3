// Josaphat Ngoga
// jngoga@g.hmc.edu
// 9/11/2025

// This module synchronizes the sequence of key inputs from the keypad and send them
// to the dual 7-segment display.

module synchronizer (
        input logic clk, reset,
        input logic [3:0] key,
        output logic [3:0] sw1, sw2);

endmodule