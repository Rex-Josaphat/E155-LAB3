// Josaphat Ngoga
// jngoga@g.hmc.edu
// 9/5/2025

